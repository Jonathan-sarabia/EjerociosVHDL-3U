
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity cont8bits_selector is
end cont8bits_selector;

architecture Behavioral of cont8bits_selector is

begin


end Behavioral;

